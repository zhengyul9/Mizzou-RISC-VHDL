    Mac OS X            	   2       9                                      ATTR      9   �   }                  �   *  com.apple.quarantine    �   S  com.dropbox.attributes   q/0082;58aa0c77;RAR\x20Extractor\x20Free; x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%G��¢(��"��˴�p�좰�@[[���Z �k�